module not_gate(output out, input in);
  nand(out, in, in);
endmodule
